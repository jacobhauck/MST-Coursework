State|Population (2016)|Population (2017)
Alabama|4860545|4874747
Alaska|741522|739795
Arizona|6908642|7016270
Arkansas|2988231|3004279
California|39296476|39536653
Colorado|5530105|5607154
Connecticut|3587685|3588184
Delaware|952698|961939
District of Columbia|684336|693972
Florida|20656589|20984400
Georgia|10313620|10429379
Hawaii|1428683|1427538
Idaho|1680026|1716943
Illinois|12835726|12802023
Indiana|6634007|6666818
Iowa|3130869|3145711
Kansas|2907731|2913123
Kentucky|4436113|4454189
Louisiana|4686157|4684333
Maine|1330232|1335907
Maryland|6024752|6052177
Massachusetts|6823721|6859819
Michigan|9933445|9962311
Minnesota|5525050|5576606
Mississippi|2985415|2984100
Missouri|6091176|6113532
Montana|1038656|1050493
Nebraska|1907603|1920076
Nevada|2939254|2998039
New Hampshire|1335015|1342795
New Jersey|8978416|9005644
New Mexico|2085432|2088070
New York|19836286|19849399
North Carolina|10156689|10273419
North Dakota|755548|755393
Ohio|11622554|11658609
Oklahoma|3921207|3930864
Oregon|4085989|4142776
Pennsylvania|12787085|12805537
Rhode Island|1057566|1059639
South Carolina|4959822|5024369
South Dakota|861542|869666
Tennessee|6649404|6715984
Texas|27904862|28304596
Utah|3044321|3101833
Vermont|623354|623657
Virginia|8414380|8470020
Washington|7280934|7405743
West Virginia|1828637|1815857
Wisconsin|5772917|5795483
Wyoming|584910|579315
Puerto Rico|3406520|3337177
